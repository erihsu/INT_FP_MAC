`timescale 1ns/10ps
//------------------------------------------------------
// define 
//------------------------------------------------------
`define CYCLE     10

module mac_tb ;
//------------------------------------------------------
// reg && wire
//------------------------------------------------------
reg  [15:0] a ,b                       ; 
reg         clk,reset                  ;
wire [15:0] mac_out                    ;


//------------------------------------------------------
// clock generation
//------------------------------------------------------
always begin #(`CYCLE/2) clk=~clk ; end  


initial begin
	a         = 'b0 ;
	b         = 'b0 ;
	clk       = 'b0 ;
	
	@(negedge clk) reset=1'b0  ;
		#(`CYCLE*2) reset=1'b1 ;
		
	@(negedge clk) ;
		{a,b}={16'b0100000101001100,16'b1001011101100010} ;

	#100;
	$finish;
end

//------------------------------------------------------
//  generate wave
//------------------------------------------------------
initial begin
   $dumpfile("mac.vcd");
   $dumpvars;
end

//------------------------------------------------------
//  Instance sram 
//------------------------------------------------------
mac_xzy u0_mac
(.clk              ( clk       )
,.rst_n             ( reset         )
,.enable              ( 1'b1       )
,.valid        ( 1'b1 )
,.read			(1'b0)
,.mode (1'b0)
,.cfg (1'b0)
,.in_a         ( a  )
,.in_b        ( b )
,.mac_out          ( mac_out   )
);


endmodule