`include "mac_if.sv"

package mac_agent_pkg;

  import uvm_pkg::*;
  `include "macro_def.sv"
  `include "mac_tr.svh"
  `include "mac_sequencer.svh"
  `include "mac_drv.svh"
  `include "mac_mon.svh"
  `include "mac_agent.svh"
  `include "mac_sequence.svh"
  
endpackage
