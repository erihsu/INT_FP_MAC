`include "mac_agent_pkg.sv"
package seq_pkg;

import uvm_pkg::*;
import mac_agent_pkg::*;

`include "base_seq.svh"


endpackage