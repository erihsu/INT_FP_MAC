// The fp16 adder not consider overflow, underflow, rounding.

module fp16_adder(a, b, c);

    input [15:0] a,b;
    output [15:0] c;

    wire a_sign, b_sign, c_sign,a_zero,b_zero;
    wire [9:0] a_mantissa, b_mantissa;
    wire [4:0] a_exponent, b_exponent, c_exponent; 

 
//

//code 

//

endmodule